* First simulation "continuous time" (from SKY130_Track_and_Hold.ipynb)
.inc track_hold_netlist_300.spice
.option method=gear
.tran {per} {per*(nfft+3)}
.end
